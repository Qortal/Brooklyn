//-----------------------------------------------------------------------------
//     The confidential and proprietary information contained in this file may
//     only be used by a person authorised under and to the extent permitted
//     by a subsisting licensing agreement from ARM Limited or its affiliates.
//
//            (C) COPYRIGHT 2015-2020 ARM Limited or its affiliates.
//                ALL RIGHTS RESERVED
//
//     This entire notice must be reproduced on all copies of this file
//     and copies of this file may only be made by a person if such person is
//     permitted to do so under the terms of a subsisting license agreement
//     from ARM Limited or its affiliates.
//
//     Release Information : HERCULESAE-MP106-r0p1-00eac0
//
//-----------------------------------------------------------------------------
// SystemVerilog (IEEE Std 1800-2012)
//-----------------------------------------------------------------------------




`include "herculesae_header.sv"


module herculesae_vx_aesimc
(


  input wire [127:0]    d_in,

  output wire [127:0]   imc 
);







  wire [7:0]                             i00;
  wire [7:0]                             i01;
  wire [7:0]                             i02;
  wire [7:0]                             i03;
  wire [7:0]                             i10;
  wire [7:0]                             i11;
  wire [7:0]                             i12;
  wire [7:0]                             i13;
  wire [7:0]                             i20;
  wire [7:0]                             i21;
  wire [7:0]                             i22;
  wire [7:0]                             i23;
  wire [7:0]                             i30;
  wire [7:0]                             i31;
  wire [7:0]                             i32;
  wire [7:0]                             i33;
  wire [7:0]                             s00;
  wire [10:0]                            s00_nr;
  wire [7:0]                             s01;
  wire [10:0]                            s01_nr;
  wire [7:0]                             s02;
  wire [10:0]                            s02_nr;
  wire [7:0]                             s03;
  wire [10:0]                            s03_nr;
  wire [7:0]                             s10;
  wire [10:0]                            s10_nr;
  wire [7:0]                             s11;
  wire [10:0]                            s11_nr;
  wire [7:0]                             s12;
  wire [10:0]                            s12_nr;
  wire [7:0]                             s13;
  wire [10:0]                            s13_nr;
  wire [7:0]                             s20;
  wire [10:0]                            s20_nr;
  wire [7:0]                             s21;
  wire [10:0]                            s21_nr;
  wire [7:0]                             s22;
  wire [10:0]                            s22_nr;
  wire [7:0]                             s23;
  wire [10:0]                            s23_nr;
  wire [7:0]                             s30;
  wire [10:0]                            s30_nr;
  wire [7:0]                             s31;
  wire [10:0]                            s31_nr;
  wire [7:0]                             s32;
  wire [10:0]                            s32_nr;
  wire [7:0]                             s33;
  wire [10:0]                            s33_nr;


assign i33[7:0] = d_in[127:120];
assign i23[7:0] = d_in[119:112];
assign i13[7:0] = d_in[111:104];
assign i03[7:0] = d_in[103:96];

assign i32[7:0] = d_in[95:88];
assign i22[7:0] = d_in[87:80];
assign i12[7:0] = d_in[79:72];
assign i02[7:0] = d_in[71:64];

assign i31[7:0] = d_in[63:56];
assign i21[7:0] = d_in[55:48];
assign i11[7:0] = d_in[47:40];
assign i01[7:0] = d_in[39:32];

assign i30[7:0] = d_in[31:24];
assign i20[7:0] = d_in[23:16];
assign i10[7:0] = d_in[15:8];
assign i00[7:0] = d_in[7:0];



assign s00_nr[10:0] = {i00[7:0],3'b000} ^ {1'b0,i00[7:0],2'b00} ^ {2'b00,i00[7:0],1'b0} 
                    ^ {i10[7:0],3'b000}                         ^ {2'b00,i10[7:0],1'b0} ^ {3'b000,i10[7:0]}
                    ^ {i20[7:0],3'b000} ^ {1'b0,i20[7:0],2'b00}                         ^ {3'b000,i20[7:0]} 
                    ^ {i30[7:0],3'b000}                                                 ^ {3'b000,i30[7:0]};
assign s00[7:0] = s00_nr[7:0] ^ ({8{s00_nr[8]}} & 8'h1b) ^ ({8{s00_nr[9]}} & 8'h36) ^ ({8{s00_nr[10]}} & 8'h6c);

assign s01_nr[10:0] = {i01[7:0],3'b000} ^ {1'b0,i01[7:0],2'b00} ^ {2'b00,i01[7:0],1'b0} 
                    ^ {i11[7:0],3'b000}                         ^ {2'b00,i11[7:0],1'b0} ^ {3'b000,i11[7:0]}
                    ^ {i21[7:0],3'b000} ^ {1'b0,i21[7:0],2'b00}                         ^ {3'b000,i21[7:0]} 
                    ^ {i31[7:0],3'b000}                                                 ^ {3'b000,i31[7:0]};
assign s01[7:0] = s01_nr[7:0] ^ ({8{s01_nr[8]}} & 8'h1b) ^ ({8{s01_nr[9]}} & 8'h36) ^ ({8{s01_nr[10]}} & 8'h6c);

assign s02_nr[10:0] = {i02[7:0],3'b000} ^ {1'b0,i02[7:0],2'b00} ^ {2'b00,i02[7:0],1'b0} 
                    ^ {i12[7:0],3'b000}                         ^ {2'b00,i12[7:0],1'b0} ^ {3'b000,i12[7:0]}
                    ^ {i22[7:0],3'b000} ^ {1'b0,i22[7:0],2'b00}                         ^ {3'b000,i22[7:0]} 
                    ^ {i32[7:0],3'b000}                                                 ^ {3'b000,i32[7:0]};
assign s02[7:0] = s02_nr[7:0] ^ ({8{s02_nr[8]}} & 8'h1b) ^ ({8{s02_nr[9]}} & 8'h36) ^ ({8{s02_nr[10]}} & 8'h6c);

assign s03_nr[10:0] = {i03[7:0],3'b000} ^ {1'b0,i03[7:0],2'b00} ^ {2'b00,i03[7:0],1'b0} 
                    ^ {i13[7:0],3'b000}                         ^ {2'b00,i13[7:0],1'b0} ^ {3'b000,i13[7:0]}
                    ^ {i23[7:0],3'b000} ^ {1'b0,i23[7:0],2'b00}                         ^ {3'b000,i23[7:0]} 
                    ^ {i33[7:0],3'b000}                                                 ^ {3'b000,i33[7:0]};
assign s03[7:0] = s03_nr[7:0] ^ ({8{s03_nr[8]}} & 8'h1b) ^ ({8{s03_nr[9]}} & 8'h36) ^ ({8{s03_nr[10]}} & 8'h6c);

assign s10_nr[10:0] = {i10[7:0],3'b000} ^ {1'b0,i10[7:0],2'b00} ^ {2'b00,i10[7:0],1'b0} 
                    ^ {i20[7:0],3'b000}                         ^ {2'b00,i20[7:0],1'b0} ^ {3'b000,i20[7:0]}
                    ^ {i30[7:0],3'b000} ^ {1'b0,i30[7:0],2'b00}                         ^ {3'b000,i30[7:0]} 
                    ^ {i00[7:0],3'b000}                                                 ^ {3'b000,i00[7:0]};
assign s10[7:0] = s10_nr[7:0] ^ ({8{s10_nr[8]}} & 8'h1b) ^ ({8{s10_nr[9]}} & 8'h36) ^ ({8{s10_nr[10]}} & 8'h6c);

assign s11_nr[10:0] = {i11[7:0],3'b000} ^ {1'b0,i11[7:0],2'b00} ^ {2'b00,i11[7:0],1'b0} 
                    ^ {i21[7:0],3'b000}                         ^ {2'b00,i21[7:0],1'b0} ^ {3'b000,i21[7:0]}
                    ^ {i31[7:0],3'b000} ^ {1'b0,i31[7:0],2'b00}                         ^ {3'b000,i31[7:0]} 
                    ^ {i01[7:0],3'b000}                                                 ^ {3'b000,i01[7:0]};
assign s11[7:0] = s11_nr[7:0] ^ ({8{s11_nr[8]}} & 8'h1b) ^ ({8{s11_nr[9]}} & 8'h36) ^ ({8{s11_nr[10]}} & 8'h6c);

assign s12_nr[10:0] = {i12[7:0],3'b000} ^ {1'b0,i12[7:0],2'b00} ^ {2'b00,i12[7:0],1'b0} 
                    ^ {i22[7:0],3'b000}                         ^ {2'b00,i22[7:0],1'b0} ^ {3'b000,i22[7:0]}
                    ^ {i32[7:0],3'b000} ^ {1'b0,i32[7:0],2'b00}                         ^ {3'b000,i32[7:0]} 
                    ^ {i02[7:0],3'b000}                                                 ^ {3'b000,i02[7:0]};
assign s12[7:0] = s12_nr[7:0] ^ ({8{s12_nr[8]}} & 8'h1b) ^ ({8{s12_nr[9]}} & 8'h36) ^ ({8{s12_nr[10]}} & 8'h6c);

assign s13_nr[10:0] = {i13[7:0],3'b000} ^ {1'b0,i13[7:0],2'b00} ^ {2'b00,i13[7:0],1'b0} 
                    ^ {i23[7:0],3'b000}                         ^ {2'b00,i23[7:0],1'b0} ^ {3'b000,i23[7:0]}
                    ^ {i33[7:0],3'b000} ^ {1'b0,i33[7:0],2'b00}                         ^ {3'b000,i33[7:0]} 
                    ^ {i03[7:0],3'b000}                                                 ^ {3'b000,i03[7:0]};
assign s13[7:0] = s13_nr[7:0] ^ ({8{s13_nr[8]}} & 8'h1b) ^ ({8{s13_nr[9]}} & 8'h36) ^ ({8{s13_nr[10]}} & 8'h6c);

assign s20_nr[10:0] = {i20[7:0],3'b000} ^ {1'b0,i20[7:0],2'b00} ^ {2'b00,i20[7:0],1'b0} 
                    ^ {i30[7:0],3'b000}                         ^ {2'b00,i30[7:0],1'b0} ^ {3'b000,i30[7:0]}
                    ^ {i00[7:0],3'b000} ^ {1'b0,i00[7:0],2'b00}                         ^ {3'b000,i00[7:0]} 
                    ^ {i10[7:0],3'b000}                                                 ^ {3'b000,i10[7:0]};
assign s20[7:0] = s20_nr[7:0] ^ ({8{s20_nr[8]}} & 8'h1b) ^ ({8{s20_nr[9]}} & 8'h36) ^ ({8{s20_nr[10]}} & 8'h6c);

assign s21_nr[10:0] = {i21[7:0],3'b000} ^ {1'b0,i21[7:0],2'b00} ^ {2'b00,i21[7:0],1'b0} 
                    ^ {i31[7:0],3'b000}                         ^ {2'b00,i31[7:0],1'b0} ^ {3'b000,i31[7:0]}
                    ^ {i01[7:0],3'b000} ^ {1'b0,i01[7:0],2'b00}                         ^ {3'b000,i01[7:0]} 
                    ^ {i11[7:0],3'b000}                                                 ^ {3'b000,i11[7:0]};
assign s21[7:0] = s21_nr[7:0] ^ ({8{s21_nr[8]}} & 8'h1b) ^ ({8{s21_nr[9]}} & 8'h36) ^ ({8{s21_nr[10]}} & 8'h6c);

assign s22_nr[10:0] = {i22[7:0],3'b000} ^ {1'b0,i22[7:0],2'b00} ^ {2'b00,i22[7:0],1'b0} 
                    ^ {i32[7:0],3'b000}                         ^ {2'b00,i32[7:0],1'b0} ^ {3'b000,i32[7:0]}
                    ^ {i02[7:0],3'b000} ^ {1'b0,i02[7:0],2'b00}                         ^ {3'b000,i02[7:0]} 
                    ^ {i12[7:0],3'b000}                                                 ^ {3'b000,i12[7:0]};
assign s22[7:0] = s22_nr[7:0] ^ ({8{s22_nr[8]}} & 8'h1b) ^ ({8{s22_nr[9]}} & 8'h36) ^ ({8{s22_nr[10]}} & 8'h6c);

assign s23_nr[10:0] = {i23[7:0],3'b000} ^ {1'b0,i23[7:0],2'b00} ^ {2'b00,i23[7:0],1'b0} 
                    ^ {i33[7:0],3'b000}                         ^ {2'b00,i33[7:0],1'b0} ^ {3'b000,i33[7:0]}
                    ^ {i03[7:0],3'b000} ^ {1'b0,i03[7:0],2'b00}                         ^ {3'b000,i03[7:0]} 
                    ^ {i13[7:0],3'b000}                                                 ^ {3'b000,i13[7:0]};
assign s23[7:0] = s23_nr[7:0] ^ ({8{s23_nr[8]}} & 8'h1b) ^ ({8{s23_nr[9]}} & 8'h36) ^ ({8{s23_nr[10]}} & 8'h6c);

assign s30_nr[10:0] = {i30[7:0],3'b000} ^ {1'b0,i30[7:0],2'b00} ^ {2'b00,i30[7:0],1'b0} 
                    ^ {i00[7:0],3'b000}                         ^ {2'b00,i00[7:0],1'b0} ^ {3'b000,i00[7:0]}
                    ^ {i10[7:0],3'b000} ^ {1'b0,i10[7:0],2'b00}                         ^ {3'b000,i10[7:0]} 
                    ^ {i20[7:0],3'b000}                                                 ^ {3'b000,i20[7:0]};
assign s30[7:0] = s30_nr[7:0] ^ ({8{s30_nr[8]}} & 8'h1b) ^ ({8{s30_nr[9]}} & 8'h36) ^ ({8{s30_nr[10]}} & 8'h6c);

assign s31_nr[10:0] = {i31[7:0],3'b000} ^ {1'b0,i31[7:0],2'b00} ^ {2'b00,i31[7:0],1'b0} 
                    ^ {i01[7:0],3'b000}                         ^ {2'b00,i01[7:0],1'b0} ^ {3'b000,i01[7:0]}
                    ^ {i11[7:0],3'b000} ^ {1'b0,i11[7:0],2'b00}                         ^ {3'b000,i11[7:0]} 
                    ^ {i21[7:0],3'b000}                                                 ^ {3'b000,i21[7:0]};
assign s31[7:0] = s31_nr[7:0] ^ ({8{s31_nr[8]}} & 8'h1b) ^ ({8{s31_nr[9]}} & 8'h36) ^ ({8{s31_nr[10]}} & 8'h6c);

assign s32_nr[10:0] = {i32[7:0],3'b000} ^ {1'b0,i32[7:0],2'b00} ^ {2'b00,i32[7:0],1'b0} 
                    ^ {i02[7:0],3'b000}                         ^ {2'b00,i02[7:0],1'b0} ^ {3'b000,i02[7:0]}
                    ^ {i12[7:0],3'b000} ^ {1'b0,i12[7:0],2'b00}                         ^ {3'b000,i12[7:0]} 
                    ^ {i22[7:0],3'b000}                                                 ^ {3'b000,i22[7:0]};
assign s32[7:0] = s32_nr[7:0] ^ ({8{s32_nr[8]}} & 8'h1b) ^ ({8{s32_nr[9]}} & 8'h36) ^ ({8{s32_nr[10]}} & 8'h6c);

assign s33_nr[10:0] = {i33[7:0],3'b000} ^ {1'b0,i33[7:0],2'b00} ^ {2'b00,i33[7:0],1'b0} 
                    ^ {i03[7:0],3'b000}                         ^ {2'b00,i03[7:0],1'b0} ^ {3'b000,i03[7:0]}
                    ^ {i13[7:0],3'b000} ^ {1'b0,i13[7:0],2'b00}                         ^ {3'b000,i13[7:0]} 
                    ^ {i23[7:0],3'b000}                                                 ^ {3'b000,i23[7:0]};
assign s33[7:0] = s33_nr[7:0] ^ ({8{s33_nr[8]}} & 8'h1b) ^ ({8{s33_nr[9]}} & 8'h36) ^ ({8{s33_nr[10]}} & 8'h6c);

assign imc[127:120] = s33[7:0];
assign imc[119:112] = s23[7:0];
assign imc[111:104] = s13[7:0];
assign imc[103:96]  = s03[7:0];

assign imc[95:88]   = s32[7:0];
assign imc[87:80]   = s22[7:0];
assign imc[79:72]   = s12[7:0];
assign imc[71:64]   = s02[7:0];

assign imc[63:56]   = s31[7:0];
assign imc[55:48]   = s21[7:0];
assign imc[47:40]   = s11[7:0];
assign imc[39:32]   = s01[7:0];

assign imc[31:24]   = s30[7:0];
assign imc[23:16]   = s20[7:0];
assign imc[15:8]    = s10[7:0];
assign imc[7:0]     = s00[7:0];

endmodule


`define HERCULESAE_UNDEFINE
`include "herculesae_header.sv"
`undef HERCULESAE_UNDEFINE
